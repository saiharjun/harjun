*** SPICE deck for cell NAND2{lay} from library Tut1
*** Created on Sat Sep 12, 2020 19:00:01
*** Last revised on Sun Sep 13, 2020 19:25:22
*** Written on Sun Sep 13, 2020 20:37:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND2{lay}
Mnmos@5 net@16 B gnd gnd nMOS L=0.4U W=2.4U AS=7.92P AD=1.2P PS=19U PD=3.4U
Mnmos@6 A_NAND_B A net@16 gnd nMOS L=0.4U W=2.4U AS=1.2P AD=2.32P PS=3.4U PD=5.133U
Mpmos@3 A_NAND_B B vdd vdd pMOS L=0.4U W=2.4U AS=5.52P AD=2.32P PS=13.2U PD=5.133U
Mpmos@4 vdd A A_NAND_B vdd pMOS L=0.4U W=2.4U AS=2.32P AD=5.52P PS=5.133U PD=13.2U

* Spice Code nodes in cell cell 'NAND2{lay}'
vdd VDD 0 DC 5 
vin A 0 pulse(0 5 10n 0.5n 0.5n 20n)
vin2 B 0 DC 5 
cload A_NAND_B 0 500ff 
.tran 0 40n 
.include c5_modeles.txt
.END
